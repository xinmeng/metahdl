module moda (
  i1, 
  i2, 
  o1, 
  o2);


input             i1;
input             i2;
output            o1;
output  [1   :0]  o2;

wire              i1;
wire              i2;
wire              o1;
wire    [1   :0]  o2;

endmodule
