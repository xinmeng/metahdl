`ifndef __xregister_vh__
`define __xregister_vh__

`define SW_RO    4'd0
`define SW_RW    4'd1
`define SW_RW1C  4'd2
`define SW_RW1S  4'd3
`define SW_ROC   4'd4
`define SW_ConC  4'd5
`define SW_WonC  4'd6

`define HW_RO     4'd0
`define HW_WIRED  4'd1
`define HW_SET    4'd2
`define HW_CLR    4'd3
`define HW_INC    4'd4
`define HW_DEC    4'd5
`define HW_ADD    4'd6
`define HW_SUB    4'd7
`define HW_VALUE  4'd8

`define SW 0
`define HW 1

`define DEBUG 1


`endif
